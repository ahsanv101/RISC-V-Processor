module registerFile
(
	input [63:0] WriteData,
	input [4:0] RS1 ,
	input [4:0] RS2,
	input [4:0] RD,
	input clk,
	input reset,
	input RegWrite,
	output reg [63:0] ReadData1,
	output reg [63:0] ReadData2

);
	reg [63:0] Register[17:0];
	initial
		begin 
			Register[0] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
			Register[1] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000001;
			Register[2] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000010;
			Register[3] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000011;
			Register[4] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000100;
			Register[5] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000101;
			Register[6] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000110;
			Register[7] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000111;
			Register[8] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001000;
			Register[9] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001001;
			Register[10] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001010;
			Register[11] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001011;
			Register[12] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001100;
			Register[13] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001101;
			Register[14] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001110;
			Register[15] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00001111;
			Register[16] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00010000;
			Register[17] = 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00010001;		
		end
always @ (posedge reset or negedge clk or RegWrite)
begin 
	if (RegWrite)
		begin
			Register[RD] = WriteData;
			ReadData1=Register[RD];
		end
	else if(!RegWrite) 
		begin
			ReadData1 = Register[RS1];
			ReadData2 =  Register[RS2];
		end
	else 
		begin
			ReadData1= 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
			ReadData2= 64'b00000000_00000000_00000000_00000000_00000000_00000000_00000000_00000000;
		end
end

endmodule